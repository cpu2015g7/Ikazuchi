library ieee;
use ieee.std_logic_1164.all;

use work.types.all;

package data is
	constant test_prog1 : rom_t := (
		"00110000000000010000000000001001",
		"00110000000000100000000000100110",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000001000100001000000100000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"11111100000000010000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		others => (others => '0')
	);

	constant loop_easy : rom_t := (
		x"3002000A",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210001",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10410004",
		x"00000000",
		x"00000000",
		x"1000FFF6",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210000",
		x"00000000",
		x"1000FFFB",
		x"00000000",
		x"00000000",
		x"00000000",
		others => (others => '0')
	);

	constant loop_hard : rom_t := (
		x"3002000A",
		x"30210001",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10410002",
		x"00000000",
		x"00000000",
		x"1000FFF7",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210000",
		x"00000000",
		x"1000FFFC",
		x"00000000",
		x"00000000",
		x"00000000",
		x"1000FFEC",
		others => (others => '0')
);

	constant fib_loop : rom_t := (
		x"3005000A",
		x"30040000",
		x"30010000",
		x"30020001",
		x"00000000",
		x"10A40006",
		x"30840001",
		x"00000000",
		x"00221820",
		x"00000000",
		x"1000FFF9",
		x"30410000",
		x"30620000",
		x"FC200000",
		x"1000FFFE",
		x"00000000",
		x"00000000",
		others => (others => '0')
);

	constant jal_test : rom_t := (
		x"3001000A",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210001",
		x"0C000001",
		others => (others => '0')
);
	constant adds_test : rom_t := (
		x"30010001",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00210820",
		x"00000000",
		x"00000000",
		x"00210820",
		x"00000000",
		x"00210820",
		x"00000000",
		x"FC200000",
		others => (others => '0')
);
	constant call_return_test : rom_t := (
		x"0C000009",
		x"00000000",
		x"00000000",
		x"00000000",
		x"1000FFFD",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10000064",
		x"30010001",
		x"00000000",
		x"00000000",
		x"03E00008",
		x"10000064",
		others => (others => '0')
);
	constant beq_test : rom_t := (
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"1000FFFD",
		x"30010001",
		x"30020001",
		x"00000000",
		others => (others => '0')
);

	constant fib_loop10_new : rom_t := (
		x"3005000A",
		x"30040000",
		x"30010000",
		x"30020001",
		x"10A40004",
		x"30840001",
		x"00221820",
		x"30410000",
		x"1000FFFA",
		x"30620000",
		x"FC200000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210001",
		x"1000FFFC",
		others => (others => '0')
);

	constant test_prog2 : rom_t := (
		x"3005000A",
		x"30040000",
		x"30010000",
		x"30020001",
		x"10A40005",
		x"30840001",
		x"00221820",
		x"30410000",
		x"1000FFFB",
		x"30620000",
		x"FC200000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210001",
		x"1000FFFF",
		others => (others => '0')
);

	constant lwsw : rom_t := (
		x"3001001E",
		x"00000000",
		x"AC010000",
		x"8C020000",
		x"8C030000",
		x"8C040000",
		x"8C050000",
		x"8C060000",
		others => (others => '0')
);
constant lwsw2 : rom_t := (
x"3009003F",
x"30010001",
x"30020002",
x"30030003",
x"AD210000",
x"AD220004",
x"AD230008",
x"8D240000",
x"8D250004",
x"8D260008",
x"00000008",
others => (others => '0')
);
	constant fib_rec : rom_t := (
x"30090200",
x"3001000A",
x"0C000007",
x"FC200000",
x"1000FFFF",
x"00000000",
x"00000000",
x"3129FFE8",
x"00000000",
x"AD3F0000",
x"AD210004",
x"10010017",
x"3021FFFF",
x"00000000",
x"00000000",
x"00000000",
x"10010012",
x"00000000",
x"0C000007",
x"00000000",
x"AD210008",
x"8D210004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3021FFFE",
x"0C000007",
x"8D220008",
x"8D3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00220820",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"31290018",
x"03E00008",

		others => (others => '0')
);

constant fib_rec2 : rom_t := (
x"30090200",
x"3001000A",
x"301D0001",
x"0C000008",
x"FC200000",
x"1000FFFF",
x"00000000",
x"00000000",
x"3129FFE8",
x"03A1182A",
x"AD3F0000",
x"AD210004",
x"10030017",
x"00000000",
x"3021FFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"0C000008",
x"00000000",
x"AD210008",
x"8D210004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3021FFFE",
x"0C000008",
x"8D220008",
x"8D3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00220820",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"31290018",
x"03E00008",
others => (others => '0')
);

end package;
