library ieee;
use ieee.std_logic_1164.all;

use work.types.all;

package data is
	constant test_prog1 : rom_t := (
		"00110000000000010000000000001001",
		"00110000000000100000000000100110",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000001000100001000000100000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"11111100000000010000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		others => (others => '0')
	);

	constant loop_easy : rom_t := (
		x"3002000A",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210001",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10410004",
		x"00000000",
		x"00000000",
		x"1000FFF6",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210000",
		x"00000000",
		x"1000FFFB",
		x"00000000",
		x"00000000",
		x"00000000",
		others => (others => '0')
	);

	constant loop_hard : rom_t := (
		x"3002000A",
		x"30210001",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10410002",
		x"00000000",
		x"00000000",
		x"1000FFF7",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210000",
		x"00000000",
		x"1000FFFC",
		x"00000000",
		x"00000000",
		x"00000000",
		x"1000FFEC",
		others => (others => '0')
);

	constant fib_loop : rom_t := (
		x"3005000A",
		x"30040000",
		x"30010000",
		x"30020001",
		x"00000000",
		x"10A40006",
		x"30840001",
		x"00000000",
		x"00221820",
		x"00000000",
		x"1000FFF9",
		x"30410000",
		x"30620000",
		x"FC200000",
		x"1000FFFE",
		x"00000000",
		x"00000000",
		others => (others => '0')
);

	constant jal_test : rom_t := (
		x"3001000A",
		x"00000000",
		x"00000000",
		x"00000000",
		x"30210001",
		x"0C000001",
		others => (others => '0')
);
	constant adds_test : rom_t := (
		x"30010001",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00210820",
		x"00000000",
		x"00000000",
		x"00210820",
		x"00000000",
		x"00210820",
		x"00000000",
		x"FC200000",
		others => (others => '0')
);
	constant call_return_test : rom_t := (
		x"0C000009",
		x"00000000",
		x"00000000",
		x"00000000",
		x"1000FFFD",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10000064",
		x"30010001",
		x"00000000",
		x"00000000",
		x"03E00008",
		x"10000064",
		others => (others => '0')
);

end package;
