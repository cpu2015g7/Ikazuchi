library ieee;
use ieee.std_logic_1164.all;

use work.types.all;

package data is

constant fib_loop : rom_t := (
		x"3005000A",
		x"30040000",
		x"30010000",
		x"30020001",
		x"00000000",
		x"10A40006",
		x"30840001",
		x"00000000",
		x"00221820",
		x"00000000",
		x"1000FFF9",
		x"30410000",
		x"30620000",
		x"FC200000",
		x"1000FFFE",
		x"00000000",
		x"00000000",
		others => (others => '0')
);

constant lwsw2 : rom_t := (
		x"3009003F",
		x"30010001",
		x"30020002",
		x"30030003",
		x"AD210000",
		x"AD220004",
		x"AD230008",
		x"8D240000",
		x"8D250004",
		x"8D260008",
		x"00000008",
		others => (others => '0')
);

constant fib_rec2 : rom_t := (
		x"3009FFFF",
		x"3001001E",
		x"0C000007",
		x"FC200000",
		x"1000FFFF",
		x"00000000",
		x"00000000",
		x"3129FFF4",
		x"00000000",
		x"AD3F0000",
		x"AD210004",
		x"10010017",
		x"3021FFFF",
		x"00000000",
		x"00000000",
		x"00000000",
		x"10010012",
		x"00000000",
		x"0C000007",
		x"00000000",
		x"AD210008",
		x"8D210004",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"3021FFFE",
		x"0C000007",
		x"8D220008",
		x"8D3F0000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00220820",
		x"00000000",
		x"00000000",
		x"00000000",
		x"00000000",
		x"3129000C",
		x"03E00008",	
		others => (others => '0')
);

end package;
