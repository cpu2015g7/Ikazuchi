library ieee;
use ieee.std_logic_1164.all;

use work.types.all;

package data is

constant tttt : rom_t := (
x"30010002",
x"00000000",
x"301D00FF",
x"00000000",
x"AFA10005",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"8C020001",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"8FAB0005",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"FD600000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"1000FFFF",
others => (others => '0')
);

constant fib_hand : rom_t := (

x"300903FF",
x"00000000",
x"3001000A",
x"00000000",
x"301D0001",
x"00000000",
x"0C000011",
x"00000000",
x"FC200000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"1000FFFE",
x"00000000",
x"00000000",
x"3129FFFA",
x"00000000",
x"03A1182A",
x"00000000",
x"AD3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"AD210001",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"1003002B",
x"00000000",
x"3021FFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"0C000011",
x"00000000",
x"00000000",
x"AD210002",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"8D210001",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3021FFFE",
x"00000000",
x"0C000011",
x"00000000",
x"8D220002",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"8D3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00220820",
x"00000000",
x"00000000",
x"31290006",
x"00000000",
x"00000000",
x"03E00008",
x"00000000",
others => (others => '0')
);

constant fib_compiler : rom_t := (

x"341D1FFF",
x"00000000",
x"00000000",
x"0C000070",
x"00000000",
x"00000000",
x"1000FFFF",
x"00000000",
x"3081FFFF",
x"00000000",
x"00000000",
x"0001082A",
x"00000000",
x"00000000",
x"14010007",
x"00000000",
x"34820000",
x"00000000",
x"00000000",
x"03E00008",
x"00000000",
x"00000000",
x"3085FFFF",
x"00000000",
x"00000000",
x"AFA40000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"34A40000",
x"00000000",
x"00000000",
x"AFBFFFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"33BDFFFE",
x"00000000",
x"00000000",
x"0C000008",
x"00000000",
x"00000000",
x"33BD0002",
x"00000000",
x"00000000",
x"8FBFFFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"34440000",
x"00000000",
x"00000000",
x"8FA50000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"30A5FFFE",
x"00000000",
x"00000000",
x"AFA4FFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"34A40000",
x"00000000",
x"00000000",
x"AFBFFFFE",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"33BDFFFD",
x"00000000",
x"00000000",
x"0C000008",
x"00000000",
x"00000000",
x"33BD0003",
x"00000000",
x"00000000",
x"8FBFFFFE",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"34440000",
x"00000000",
x"00000000",
x"8FA5FFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00A41020",
x"00000000",
x"00000000",
x"03E00008",
x"00000000",
x"00000000",
x"3004000A",
x"00000000",
x"00000000",
x"AFBF0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"33BDFFFF",
x"00000000",
x"00000000",
x"0C000008",
x"00000000",
x"00000000",
x"33BD0001",
x"00000000",
x"00000000",
x"8FBF0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"34440000",
x"00000000",
x"00000000",
x"AFBF0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"33BDFFFF",
x"00000000",
x"00000000",
x"FC800000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"33BD0001",
x"00000000",
x"00000000",
x"8FBF0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"03E00008",
x"00000000",
x"00000000",
others => (others => '0')
);

constant plusone : rom_t := (
x"0C000008",
x"00000000",
x"30840064",
x"00000000",
x"3082FF9D",
x"00000000",
x"03E00008",
x"00000000",
x"3004000A",
x"00000000",
x"AFBF0004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"0C000002",
x"00000000",
x"33BD0008",
x"00000000",
x"33BDFFFF",
x"00000000",
x"8FBF0004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"34440000",
x"00000000",
x"AFBF0004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"FC800000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"33BD0008",
x"00000000",
x"33BDFFFF",
x"00000000",
x"8FBF0004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"1000FFFF",
x"00000000",
x"03E00008",
x"00000000",
others => (others => '0')
);

constant loop_back : rom_t := (
x"F8010000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"FC200000",
x"1000FFF9",
others => (others => '0')
);

constant float_io : rom_t := (

x"0C000007",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"1000FFFA",
x"00000000",
x"00000000",
x"00000000",
x"AC1F0000",
x"0C00005B",
x"00000000",
x"00000000",
x"0C00004B",
x"00000000",
x"00000000",
x"30230000",
x"0C00005B",
x"00000000",
x"00000000",
x"0C00004B",
x"00000000",
x"00000000",
x"30220000",
x"30610000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"2C221820",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"2C222001",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"2C222803",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"2C223018",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"2C223808",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"30610000",
x"0C00004B",
x"30810000",
x"0C00004B",
x"30A10000",
x"0C00004B",
x"30C10000",
x"0C00004B",
x"30E10000",
x"0C00004B",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"8C1F0000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"03E00008",
x"00000000",
x"0001D602",
x"0001CC02",
x"0001C202",
x"0001B802",
x"00000000",
x"00000000",
x"00000000",
x"FF400000",
x"FF200000",
x"FF000000",
x"FEE00000",
x"00000000",
x"00000000",
x"00000000",
x"03E00008",
x"00000000",
x"00000000",
x"F8010000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00010A00",
x"00000000",
x"F8010000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00010A00",
x"00000000",
x"F8010000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00010A00",
x"00000000",
x"F8010000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"03E00008",
others => (others => '0')
);

constant float_test : rom_t := (

x"3401D8EF",
x"34020002",
x"00010C00",
x"00021400",
x"34210014",
x"3442000F",
x"340303FF",
x"00000000",
x"00000000",
x"0C000016",
x"00000000",
x"2C221801",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"30610000",
x"00000000",
x"0C000016",
x"00000000",
x"00000000",
x"1000FFFE",
x"00000000",
x"0001D602",
x"0001CC02",
x"0001C202",
x"0001B802",
x"00000000",
x"00000000",
x"00000000",
x"FF400000",
x"FF200000",
x"FF000000",
x"FEE00000",
x"00000000",
x"00000000",
x"00000000",
x"03E00008",
others => (others => '0')
);
constant fadd_test : rom_t := (

x"3401D8EF",
x"34020002",
x"00010C00",
x"00021400",
x"34210014",
x"3442000F",
x"00000000",
x"00000000",
x"2C221808",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00032202",
x"00032C02",
x"00033602",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"FCC00000",
x"FCA00000",
x"FC800000",
x"FC600000",
x"00000000",
x"1000FFFE",
others => (others => '0')
);

constant shift_test : rom_t := (
x"30010005",
x"30020014",
x"00000000",
x"00000000",
x"00010880",
x"00021082",
x"00000000",
x"00000000",
x"00000000",
x"FC200000",
x"00000000",
x"00000000",
x"1000FFFE",
others => (others => '0')
);
constant fib_loop : rom_t := (
		x"3005000A",
		x"30040000",
		x"30010000",
		x"30020001",
		x"00000000",
		x"10A40006",
		x"30840001",
		x"00000000",
		x"00221820",
		x"00000000",
		x"1000FFF9",
		x"30410000",
		x"30620000",
		x"FC200000",
		x"1000FFFE",
		x"00000000",
		x"00000000",
		others => (others => '0')
);

constant lwsw2 : rom_t := (
		x"3009003F",
		x"30010001",
		x"30020002",
		x"30030003",
		x"AD210000",
		x"AD220004",
		x"AD230008",
		x"8D240000",
		x"8D250004",
		x"8D260008",
		x"00000008",
		others => (others => '0')
);

constant fib_rec2 : rom_t := (

x"3009FFFF",
x"3001000A",
x"0C000007",
x"FC200000",
x"FC200000",
x"1000FFFF",
x"00000000",
x"00000000",
x"3129FFF4",
x"00000000",
x"AD3F0000",
x"AD210004",
x"10010017",
x"3021FFFF",
x"00000000",
x"00000000",
x"00000000",
x"10010012",
x"00000000",
x"0C000007",
x"00000000",
x"AD210008",
x"8D210004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3021FFFE",
x"0C000007",
x"8D220008",
x"8D3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00220820",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3129000C",
x"03E00008",
		others => (others => '0')
);

constant fib_rec_old : rom_t := (

x"30097FF8",
x"30010020",
x"301D0001",
x"0C000008",
x"FC200000",
x"FC200000",
x"1000FFFF",
x"00000000",
x"00000000",
x"3129FFE8",
x"03A1182A",
x"AD3F0000",
x"AD210004",
x"10030017",
x"00000000",
x"3021FFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"0C000008",
x"00000000",
x"AD210008",
x"8D210004",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3021FFFE",
x"0C000008",
x"8D220008",
x"8D3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00220820",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"31290018",
x"03E00008",

others => (others => '0')
);

constant fib_b : rom_t := (

x"30097FF8",
x"3001001E",
x"301D0001",
x"0C000008",
x"FC200000",
x"1000FFFF",
x"00000000",
x"00000000",
x"3129FFFD",
x"03A1182A",
x"AD3F0000",
x"AD210001",
x"10030017",
x"00000000",
x"3021FFFF",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"0C000008",
x"00000000",
x"AD210002",
x"8D210001",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"3021FFFE",
x"0C000008",
x"8D220002",
x"8D3F0000",
x"00000000",
x"00000000",
x"00000000",
x"00220820",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"31290003",
x"03E00008",
others => (others => '0')
);

constant rx_tx : rom_t := (
x"30030001",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"F8030000",
x"00000000",
x"00000000",
x"FC600000",
x"1000FFFA",
others => (others => '0')
);

end package;
